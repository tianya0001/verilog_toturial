module eeprom (
    input wire sys_clk,
    input wire sys_rst,
    
    inout reg sda,
    output reg scl
);
    

    
endmodule //eeprom



